// File        :mailbox.sv
// Author      :Roopashri.C /1BM23EC218
// Created     :02-02-2026
// Module      :mailbox
// Project     :SystemVerilog & Verification(23EC6PE2SV)
// Faculty     :Prof.Ajaykumar Devarapalli
// Description :Packet class models randomized transaction data used for communication.
class Packet;
  rand bit [7:0] val;
endclass


 
